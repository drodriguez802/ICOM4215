module ram_256 (output reg[31:0] DataOut,output reg MOC,input [31:0] DataIn,input R_W,input MOV,input [7:0] Address,input [1:0] size,state);
    reg[7:0] Mem[0:255];

    // For loading instructions to RAM
    integer fd, code;
    reg[7:0] data, ptr;

    // Task to print memory contents
    task print_memory;
    begin
        ptr = 0;
        $display("Address  | Content");
        $display("----------------------------------------------");
        repeat(20) begin
            $write("%d      | ", ptr);
            repeat(4) begin
                $write("%b ", Mem[ptr]);
                ptr = ptr + 1;
            end
            $write("\n");
        end
        $display("\n");
    end
    endtask

    always @(MOV, R_W)
        begin
            if (MOV)
                begin
                    if(R_W)
                    begin
                        case(size)
                            // READING
                            // Byte
                            2'b00:
                                begin
                                    //$display("STATE: %d MAR: %d DATAOUT: %b",state,Address,DataIn);
                                    DataOut[7:0] <= Mem[Address];
                                    DataOut[31:8] <= 24'b0;
                                end
                            // Halfword
                            2'b01:
                                begin
                                    DataOut[15:8] <= Mem[Address];
                                    DataOut[7:0] <= Mem[Address + 1];
                                    DataOut[31:16] <= 16'b0;
                                end
                            // Word
                            2'b10:
                                begin
                                    DataOut[31:24] <= Mem[Address];
                                    DataOut[23:16] <= Mem[Address+1];
                                    DataOut[15:8] <= Mem[Address+2];
                                    DataOut[7:0] <= Mem[Address+3];
                                end

                        endcase
                        end
                    else
                    begin
                        case(size)
                            // WRITING
                            // Byte
                            2'b00:begin
                                Mem[Address] = DataIn[7:0];
                                $display("MAR: %d DATAIN: %b    ACTUAL: %b",Address,DataIn[7:0],Mem[Address]);
                                end

                            // Halfword
                            2'b01:
                                begin
                                    Mem[Address] <= DataIn[15:8];
                                    Mem[Address + 1] <= DataIn[7:0];
                                end
                            // Word
                            2'b10:
                                begin
                                    Mem[Address] <= DataIn[31:24];
                                    Mem[Address+1] <= DataIn[23:16];
                                    Mem[Address+2] <= DataIn[15:8];
                                    Mem[Address+3] <= DataIn[7:0];
                                end
                        endcase
                        end
                    // Turn MOC on After Operation was successful
                    MOC = 1;
                end
            else
                begin
                    //DataOut = 32'bz;
                    MOC = 0;
                end

        end

    initial begin
        ptr = 0;
        // Load RAM with instructions ------------------------------------------
        fd = $fopen("testcode_arm1.txt", "r");//change here check this
        while(!($feof(fd)) && $fscanf(fd, "%b", data)) begin
            Mem[ptr] = data;
            ptr = ptr + 1;
        end

    // Print Initial Memory Contents ---------------------------------------
        $display("----------------------------------------------");
        $display("\nInitial memory content. Instructions Loaded.\n");
        print_memory();

        #100000  // Increment time delay if necessary.
        // Print Final Memory Contents -----------------------------------------
        $display("----------------------------------------------");
        $display("\nFinal memory content.\n");
        print_memory();
    end

endmodule


module arithmetic_logic_unit (output reg [31: 0] out, output reg zero, n, c, v, input [31: 0] A, B, input [4: 0] Op, input Cin);
//Setting the conditional codes to 0 initially.

//Setting interconexions
reg [31: 0] temp;
reg  signed [31: 0] pctemp;
wire [31: 0]  zero_num;
assign zero_num=32'b00000000000000000000000000000000;

always@(A,B,Op,Cin)
begin
//Case for defining the operation to be executed
case(Op)
//AND
5'b00000:
begin
out = A & B;
c = Cin;
v = 1'b0;
end

//XOR
5'b00001:
begin
out = A ^ B;
c = Cin;
v = 1'b0;
end

//Subtract
5'b00010:
begin
c = Cin;
{c, out} = A - B;
c = ~c;
if(A[31]!=B[31])
if(B[31]==out[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//Reverse Subtract
5'b00011:
begin
c = Cin;
{c, out} = B - A;
c = ~c;
if(A[31]!=B[31])
if(A[31]==out[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//ADD
5'b00100:
begin
c = Cin;
{c, out} = A + B;
if(A[31]==B[31])
if(out[31]!=B[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//ADD w/ Carry
5'b00101:
begin
c = Cin;
{c, out} = A + B + Cin;
if(A[31]==B[31])
if(out[31]!=B[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//Subtract w/ Carry
5'b00110:
begin
c = Cin;
{c, out} = A - B - !Cin;
c = ~c;
if(A[31]!=B[31])
if(B[31]==out[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//Reverse subtract w/ Carry
5'b00111:
begin
c = Cin;
{c, out} = B - A - !Cin;
c = ~c;
if(A[31]!=B[31])
if(A[31]==out[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//Test
5'b01000:
begin
temp = A & B;
c = Cin;
v = 1'b0;
end

//Test Equivalence
5'b01001:
begin
temp = A ^ B;
c = Cin;
v = 1'b0;
end

//Compare
5'b01010:
begin
c = Cin;
{c, temp} = A - B;
c = ~c;
if(A[31]!=B[31])
if(B[31]==temp[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//Compare Negated
5'b01011:
begin
c = Cin;
{c, temp} = A + B;
if(A[31]==B[31])
if(temp[31]!=B[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//OR
5'b01100:
begin
out = A | B;
c = Cin;
v = 1'b0;
end

//Move
5'b01101:
begin
out = B;
c = Cin;
v = 1'b0;
end

//Bit Clear
5'b01110:
begin
out = A & ~B;
c = Cin;
v = 1'b0;
end

//Move Not
5'b01111:
begin
out = ~B;
c = Cin;
v = 1'b0;
end

//A
5'b10000:
begin
out = A;
c = Cin;
end

//A + 4
5'b10001:
begin
{c, out} = A + 32'b00000000000000000000000000000100;
if(A[31]==B[31])
if(out[31]!=B[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//A + B + 4
5'b10010:
begin
{c, out} = A + B + 32'b00000000000000000000000000000100;
if(A[31]==B[31])
if(out[31]!=B[31])
v=1'b1;
else v=1'b0;
else v=1'b0;
end

//Signed A*4 + B (Add an offset to PC)
5'b10011:
begin
pctemp = B * 32'h4;
out = pctemp + A;
end
endcase

//Setting the condition codes:
//N
if((Op<5'b01000) || (Op>5'b01011)) n = out[31];
else n = temp[31];
//Z
// begin
zero = ~out & ~zero_num;
//     end
// else
// begin
//     zero = 0;
//     end
//$display("A: %b B: %b OUT: %b",A,B,out);
end
endmodule

module registerfile(R5,R0,R3,R2,R1,R15,R0e,R1e,portC, portA, portB, decS3, decS2, decS1, decS0, muxAS3, muxAS2, muxAS1, muxAS0, muxBS3, muxBS2, muxBS1, muxBS0, enable, clk);
  output wire [31:0] portA, portB;
  input wire decS3;
  input wire decS2;
  input wire decS1;
  input wire decS0;
  input wire muxAS3, muxAS2, muxAS1, muxAS0, muxBS3, muxBS2, muxBS1, muxBS0;
  input wire clk, enable;
  input wire [31:0] portC;
  output wire [31:0]R0,R2,R3, R1,R15,R5;
  wire[31:0]  R4, R6, R7, R8, R9, R10, R11, R12, R13, R14;//Register Data
  output wire R0e, R1e;
  wire R2e, R3e, R4e, R5e, R6e, R7e, R8e, R9e, R10e, R11e, R12e, R13e, R14e, R15e;//enable for register Rn

  decoder #1registerFileDecoder(R0e, R1e, R2e, R3e, R4e, R5e, R6e, R7e, R8e, R9e, R10e, R11e, R12e, R13e, R14e, R15e, decS3, decS2, decS1, decS0, enable, clk);

  register #1register0(R0, portC, R0e, clk);
  register #1register1(R1, portC, R1e, clk);
  register #1register2(R2, portC, R2e, clk);
  register #1register3(R3, portC, R3e, clk);
  register #1register4(R4, portC, R4e, clk);
  register #1register5(R5, portC, R5e, clk);
  register #1register6(R6, portC, R6e, clk);
  register #1register7(R7, portC, R7e, clk);
  register #1register8(R8, portC, R8e, clk);
  register #1register9(R9, portC, R9e, clk);
  register #1register10(R10, portC, R10e, clk);
  register #1register11(R11, portC, R11e, clk);
  register #1register12(R12, portC, R12e, clk);
  register #1register13(R13, portC, R13e, clk);
  register #1register14(R14, portC, R14e, clk);
  register #1register15(R15, portC, R15e, clk);
  mux16x1 #1muxA(portA, R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, muxAS3, muxAS2, muxAS1, muxAS0);
  mux16x1 #1muxB(portB, R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, muxBS3, muxBS2, muxBS1, muxBS0);
  endmodule


module decoder(R0e, R1e, R2e, R3e, R4e, R5e, R6e, R7e, R8e, R9e, R10e, R11e, R12e, R13e, R14e, R15e, S3, S2, S1, S0, enable, clk);
        input wire S3, S2, S1, S0, enable, clk;
        output wire R0e, R1e, R2e, R3e, R4e, R5e, R6e, R7e, R8e, R9e, R10e, R11e, R12e, R13e, R14e, R15e;

        assign R0e = enable&&~S0&&~S1&&~S2&&~S3&&1'b1;//0000 - R0
        assign R1e= enable&&S0&&~S1&&~S2&&~S3&&1'b1;//0001 - R1
        assign R2e= enable&&~S0&&S1&&~S2&&~S3&&1'b1;//0010 - R2
        assign R3e= enable&&S0&&S1&&~S2&&~S3&&1'b1;//0011 - R3
        assign R4e= enable&&~S0&&~S1&&S2&&~S3&&1'b1;//0100 - R4
        assign R5e= enable&&S0&&~S1&&S2&&~S3&&1'b1;//0101 - R5
        assign R6e= enable&&~S0&&S1&&S2&&~S3&&1'b1;//0110 - R6
        assign R7e= enable&&S0&&S1&&S2&&~S3&&1'b1;//0111 - R7
        assign R8e= enable&&~S0&&~S1&&~S2&&S3&&1'b1;//1000 - R8
        assign R9e= enable&&S0&&~S1&&~S2&&S3&&1'b1;//1001 - R9
        assign R10e= enable&&~S0&&S1&&~S2&&S3&&1'b1;//1010 - R10
        assign R11e= enable&&S0&&S1&&~S2&&S3&&1'b1;//1011 - R11
        assign R12e= enable&&~S0&&~S1&&S2&&S3&&1'b1;//1100 - R12
        assign R13e= enable&&S0&&~S1&&S2&&S3&&1'b1;//1101 - R13
        assign R14e= enable&&~S0&&S1&&S2&&S3&&1'b1;//1110 - R14
        assign R15e= enable&&S0&&S1&&S2&&S3&&1'b1;//1111 - R015


endmodule


module register(out, in, enable, clk);
   input wire [31:0] in;
   input wire enable, clk;
   output reg [31:0] out = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
   always@(posedge clk)
    begin
        if(enable==1'b1)
        begin
            //$display("REGIN: %b",in);
            out <= in;
        end
    end
endmodule

module rfmultiplexer4x1(outR, inR0, inR1, inR2, inR3, S1, S0);
   input wire S1, S0;
   input [31:0] inR0, inR1, inR2, inR3;
   output reg [31:0] outR;
   wire [1:0] select;
   assign select[0] = S0;
   assign select[1] = S1;
   always@(select or inR0 or inR1 or inR2 or inR3)
    begin
        case(select)
            2'b00 : outR = inR0;
            2'b01 : outR = inR1;
            2'b10 : outR = inR2;
            2'b11 : outR = inR3;
    endcase
    end
endmodule

module rfMux(outR, inR0, inR1, inR2, inR3, S1, S0);
   input wire S1, S0;
   input [3:0] inR0, inR1, inR2, inR3;
   output reg [3:0] outR;
   wire [1:0] select;
   assign select[0] = S0;
   assign select[1] = S1;
   always@(select or inR0 or inR1 or inR2 or inR3)
    begin
        case(select)
            2'b00 : outR = inR0;
            2'b01 : outR = inR1;
            2'b10 : outR = inR2;
            2'b11 : outR = inR3;
    endcase
    end
endmodule

module mux16x1(outR, inR0, inR1, inR2, inR3, inR4, inR5, inR6, inR7,
inR8, inR9, inR10, inR11, inR12, inR13, inR14, inR15, S3, S2, S1, S0);
   input wire S3, S2, S1, S0;
   input [31:0] inR0, inR1, inR2, inR3, inR4, inR5, inR6, inR7,
inR8, inR9, inR10, inR11, inR12, inR13, inR14, inR15;
   output wire [31:0] outR;
   wire [31:0] zero, one, two, three;
   wire [3:0] select;

   rfmultiplexer4x1 muxZero(zero, inR0, inR1, inR2, inR3, S1, S0);
   rfmultiplexer4x1 muxOne(one, inR4, inR5, inR6, inR7, S1, S0);
   rfmultiplexer4x1 muxTwo(two, inR8, inR9, inR10, inR11, S1, S0);
   rfmultiplexer4x1 muxThree(three, inR12, inR13, inR14, inR15, S1, S0);
   rfmultiplexer4x1 muxFinal(outR, zero, one, two, three, S3, S2);

endmodule

//ROM For Load immediate Offset and Register Offset
module encoder(instruction, state);
   output reg [7:0]state;
   input wire [31:0] instruction;

   always@(instruction)
    begin
        //$display("INSTRUCCION: %b",instruction);
        if(instruction[27:25]==3'b001)
            begin
            //$display("STATE 5");
            state = 8'b00000101;
            end
        else if(instruction[27:25]==3'b011)
            begin
            //$display("STATE 6");
            state = 8'b00000110;
            end
        else if(instruction[27:25]==3'b010 && instruction[20]==1'b1)
        begin
            state = 8'b00001010;
        end
        else if(instruction[27:25]==3'b010 && instruction[20]==1'b0)
        begin
            state = 8'b00010100;
        end
        else if(instruction[27:25]==3'b000)
        begin
            state = 8'b00001100;
        end
        else if(instruction[27:25]==3'b101)
        begin
            state = 8'b00001101;
        end
        //$display("STATE: %b", state);
    end
endmodule

module ROM(R15,R3,zero,DataType,currentState,MA,MB,MC,MBS,MBSMRF,MUXMDR,MDREn,MAREn,IREn,SHF_S,ShiftEn,RFEn,RW,MemEn,MOV, Inv, N2, N1, N0,SignExtSel,CR,OP, state, clk,S1,S0,instruction);
   output reg MBS = 1'b0,  MUXMDR = 0, MDREn = 0, MAREn = 0, IREn = 1'b0, Inv=1'b0, N2=0, N1=1, N0=1, S1 = 1'b0, S0 = 1'b0,ShiftEn = 0,RFEn = 1'b1,RW = 0, MemEn = 0, MOC = 1, MOV = 1;
   output reg [1:0]SignExtSel = 2'b00,MA = 2'b00, MB = 2'b10,MBSMRF = 2'b00,DataType = 2'b10;
   output reg [2:0] MC = 3'b001,SHF_S = 3'b000;
   output reg [5:0] CR = 6'b000001;
   output reg [4:0]OP = 5'b01101;
   output reg [7:0] currentState = 8'b00000000;
   input wire [7:0] state;
   input wire [31:0] instruction,R3,R15;
   input wire clk,zero;

   always@(posedge clk)
    begin
        if(state==8'b00000000)
            begin
            currentState = 8'b00000000;
            MA = 2'b00;
            MB = 2'b10;
            MC = 2'b01;
            MBS = 1'b1;
            MBSMRF = 2'b10;
            MUXMDR = 0;
            DataType = 2'b10;
            MDREn = 0;
            MAREn = 1;
            IREn = 1'b0;
            SHF_S = 3'b001;
            ShiftEn = 1'b1;
            SignExtSel = 2'b10;
            RFEn = 1'b1;
            OP = 5'b01101;
            RW = 1;
            MemEn = 0;
            MOC = 1;
            MOV = 0;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b000001;
            end
        else if(state==8'b0000001)
            begin
            currentState = 8'b00000001;
            MA = 2'b10;
            MB = 2'b00;
            MC = 2'b00;
            MBS = 1'b0;
            MBSMRF = 1'b0;
            MUXMDR = 0;
            MDREn = 0;
            MAREn = 1'b1;
            IREn = 1'b1;
            SHF_S = 3'b000;
            ShiftEn = 0;
            SignExtSel = 2'b00;
            RFEn = 1'b0;
            OP = 5'b10000;
            DataType = 2'b10;
            RW = 1'b1;
            MemEn = 0;
            MOC = 1'b1;
            MOV = 1'b1;
            N2 = 0;
            N1 = 1;
            N0 = 1;
            Inv = 0;
            S1 = 0;
            S0 = 0;
            CR = 6'b000010;
            end
        else if(state==8'b0000010)
            begin
            currentState = 8'b00000010;
            MA = 2'b10;
            MB = 2'b00;
            MC = 2'b01;
            MBS = 1'b0;
            MBSMRF = 1'b0;
            MUXMDR = 0;
            MDREn = 0;
            MAREn = 0;
            IREn = 1'b0;
            SHF_S = 3'b000;
            ShiftEn = 0;
            SignExtSel = 2'b00;
            RFEn = 1'b1;
            OP = 5'b10001;
            MemEn = 1'b0;
            N2 = 0;
            N1 = 1;
            N0 = 1;
            Inv = 0;
            S1 = 0;
            S0 = 0;
            CR = 6'b000011;
            end
        else if(state==8'b00000011)
            begin
            currentState = 8'b00000011;
            MA = 2'b00;
            MB = 2'b00;
            MC = 2'b00;
            MBS = 1'b0;
            MBSMRF = 1'b0;
            MUXMDR = 0;
            MDREn = 0;
            MAREn = 0;
            IREn = 1'b1;
            SHF_S = 3'b000;
            ShiftEn = 0;
            SignExtSel = 2'b00;
            RFEn = 1'b0;
            OP = 5'b10001;
            RW = 1;
            MemEn = 1;
            MOC = 1;
            MOV = 1;
            N2 = 0;
            N1 = 1;
            N0 = 1;
            Inv = 0;
            S1 = 0;
            S0 = 0;
            CR = 6'b000100;
            end
        else if(state==8'b00000100)
            begin
            currentState = 8'b00000100;
            MA = 2'b00;
            MB = 2'b00;
            MC = 2'b00;
            MBS = 1'b0;
            MBSMRF = 1'b0;
            MUXMDR = 0;
            MDREn = 0;
            MAREn = 0;
            IREn = 1'b1;
            SHF_S = 3'b000;
            ShiftEn = 0;
            SignExtSel = 2'b00;
            RFEn = 1'b0;
            OP = 5'b10001;
            RW = 0;
            MemEn = 0;
            MOC = 0;
            MOV = 0;
            N2 = 0;
            N1 = 0;
            N0 = 0;
            Inv = 0;
            S1 = 0;
            S0 = 1;
            CR = 6'b000001;
            end

         else if(state==8'b00000101)
            begin
            currentState = 8'b00000101;
            MA = 2'b00;
            MB = 2'b01;
            MC = 2'b00;
            MBS = 1'b1;
            MBSMRF = 2'b10;
            MUXMDR = 0;
            MDREn = 0;
            MAREn = 1'b0;
            IREn = 1'b0;
            SHF_S = 3'b001;
            ShiftEn = 1'b1;
            SignExtSel = 2'b10;
            DataType = 2'b00;
            RFEn = 1'b1;
            OP = {1'b0,instruction[24:21]};
            RW = 1;
            MemEn = 1'b0;
            MOC = 1;
            MOV = 1;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b000001;
            end
        else if(state==8'b00000110)
            begin
            currentState = 8'b00000110;
            MC = 2'b00;
            MA= 2'b00;
            MB = 2'b01;
            SHF_S = 3'b001;
            IREn = 1'b0;
            OP = 5'b00100;
            DataType = 2'b00;
            RFEn = 1'b0;
            MemEn = 1'b0;
            MAREn = 1'b1;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b00000111;
            end
        else if(state==8'b00000111)
            begin
            currentState = 8'b00000111;
            MB=2'b11;
            IREn = 1'b0;
            OP = 5'b01101;
            DataType = 2'b00;
            RFEn = 1'b1;
            RW = 1'b1;
            MemEn = 1'b1;
            MAREn = 1'b0;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b000001;
            end
        else if(state==8'b00001010)
            begin
            currentState = 8'b00001010;
            MA = 2'b00;
            MC = 2'b00;
            MB = 2'b11;
            SHF_S = 3'b011;
            IREn = 1'b0;
            OP = 5'b00100;
            DataType = 2'b00;
            RFEn = 1'b0;
            RW = instruction[20];
            MemEn = 1'b0;
            MAREn = 1'b1;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b001011;
            end
        else if(state==8'b00001011)
            begin
            currentState = 8'b00001011;
            MA = 2'b00;
            IREn = 1'b0;
            RW = instruction[20];
            OP = 5'b10000;
            RFEn = 1'b0;
            MemEn = 1'b1;
            MAREn = 1'b0;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b001111;
            end
        else if(state==8'b00001111)
            begin
            currentState = 8'b00001111;
            MA = 2'b00;
            MB = 2'b11;
            IREn = 1'b0;
            OP = 5'b01101;
            RW = instruction[20];
            RFEn = instruction[20];
            MemEn = 1'b1;
            MAREn = 1'b0;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b000001;
            end
        else if(state==8'b00001100)
            begin
            currentState = 8'b00001100;
            MA = 2'b00;
            MB = 2'b00;
            MC = 2'b00;
            MBS = 1'b1;
            MBSMRF = 2'b10;
            MUXMDR = 0;
            MDREn = 0;
            MAREn = 1'b0;
            IREn = 1'b0;
            SHF_S = 3'b011;
            ShiftEn = 1'b1;
            SignExtSel = 2'b10;
            DataType = 2'b00;
            RFEn = 1'b1;
            OP = {1'b0,instruction[24:21]};
            RW = 1;
            MemEn = 1'b0;
            MOC = 1;
            MOV = 1;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b000001;
            end
        else if(state==8'b00001101)
            begin
            //$display("ZERO: %b",zero);
            if(R3!=8'h00000000||instruction==32'b11101010111111111111111111111111)
            begin
            currentState = 8'b00001101;
            MA = 2'b00;
            MB = 2'b01;
            MC = 2'b01;
            IREn = 1'b0;
            SHF_S = 3'b100;
            ShiftEn = 1'b1;
            SignExtSel = 2'b10;
            DataType = 2'b00;
            RFEn = 1'b1;
            OP = 5'b10011;
            end
            else if(R15==32'b10001000000000000000000000101000 || R15==32'b01000100000000000000000000101000)
            begin
            //$display("ITS R15");
            MA = 2'b10;
            MC = 2'b01;
            IREn = 1'b0;
            SHF_S = 3'b100;
            ShiftEn = 1'b1;
            SignExtSel = 2'b10;
            DataType = 2'b00;
            RFEn = 1'b1;
            MAREn = 1'b0;
            OP = 5'b10001;
            end
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b000001;
            end
        else if(state==8'b00010100)
            begin
            currentState = 8'b00010100;
            MA = 2'b00;
            MC = 2'b00;
            MB = 2'b11;
            SHF_S = 3'b011;
            IREn = 1'b0;
            OP = 5'b00100;
            DataType = 2'b00;
            RFEn = 1'b0;
            RW = 1'b0;
            MemEn = 1'b0;
            MAREn = 1'b1;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b010101;
            end
        else if(state==8'b00010101)
            begin
            currentState = 8'b00010101;
            MA = 2'b01;
            IREn = 1'b0;
            OP = 5'b10000;
            RFEn = 1'b0;
            MemEn = 1'b0;
            MAREn = 1'b0;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b010110;
            end
        else if(state==8'b00010110)
            begin
            currentState = 8'b00010110;
            MemEn = 1'b1;
            MAREn = 1'b0;
            N2 = 0;
            N1 = 1;
            N0 = 0;
            Inv = 0;
            S1 = 1;
            S0 = 0;
            CR = 6'b000001;
            end
    end
endmodule

module multiplexer4x1(outR, inR0, inR1, inR2, inR3, select);
   input wire S1, S0;
   input [7:0] inR0, inR1, inR2, inR3;
   output reg [7:0] outR = 8'b00000000;
   input [1:0] select;
   always@(select or inR0 or inR1 or inR2 or inR3)
    begin
        case(select)
            2'b00 : outR = inR0;
            2'b01 : outR = inR1;
            2'b10 : outR = inR2;
            2'b11 : outR = inR3;
    endcase
     //$display("SELECT WAS: %b AND OUT WAS: %b",select, outR);
    end
endmodule

module multiplexerB(outR, inR0, inR1, inR2, inR3, select);
   input wire S1, S0;
   input [31:0] inR0, inR1, inR2, inR3;
   output reg [31:0] outR = 8'h00000000;
   input [1:0] select;
   always@(select or inR0 or inR1 or inR2 or inR3)
    begin
        case(select)
            2'b00 : outR = inR0;
            2'b01 : outR = inR1;
            2'b10 : outR = inR2;
            2'b11 : outR = inR3;
    endcase
     //$display("SELECT WAS: %b AND OUT WAS: %b",select, outR);
    end
endmodule

module adder(input [7:0] value,input [7:0] one,output  [7:0] result);
        wire [7:0]result2 = value + one;
        assign result = result2;
endmodule

//Next State Address Selector
module nextStAddSel(M, Sts, N2, N1, N0);
   input wire Sts;
   input wire S1, S0;
   input wire N2, N1, N0;
   output reg [1:0] M;
   wire [2:0] nSelect;
   assign nSelect[0] = N0;
   assign nSelect[1] = N1;
   assign nSelect[2] = N2;
   always@(nSelect or N2 or N1 or N0)
    begin
        if(nSelect==000)
            M<=00;
        else if(nSelect==3'b001)
            M<=01;
        else if(nSelect==3'b010)
            M<=10;
        else if(nSelect==3'b011)
            M=11;
        else if(nSelect==3'b100 && ~Sts)
            M=00;
        else if(nSelect==3'b100 && Sts)
            M=10;
        else if(nSelect==3'b101 && ~Sts)
            M=11;
        else if(nSelect==3'b101 && Sts)
            M=10;
        else if(nSelect==3'b110 && ~Sts)
            M=11;
        else if(nSelect==3'b110 && Sts)
            M=00;
        else if(nSelect==3'b111)
            M=00;
        //$display("NEXT ADDRESS IS: %b",M);
    end
endmodule

module inverter(iBit, inv, oBit);
    input wire iBit, inv;
    output reg oBit;
    always@(iBit or inv)
    begin
        if(inv==1'b1)
            oBit=~iBit;
        else if(inv==1'b0)
            oBit=iBit;
    //$display("INVERTER IN: %b",iBit);
    //$display("INVERTER OUT: %b",oBit);
    end
endmodule

module conditionMux(outR, inR0, inR1, inR2, inR3, select);
   input wire S1, S0;
   input inR0, inR1, inR2, inR3;
   output reg outR;
   input [1:0] select;
   always@(select or inR0 or inR1 or inR2 or inR3)
    begin
        case(select)
            2'b00 : outR = inR0;
            2'b01 : outR = inR1;
            2'b10 : outR = inR2;
            2'b11 : outR = inR3;
    endcase
     //$display("CONDITIONSELECT WAS: %b",select);
     //$display("CONDITIONMUX OUT: %b",outR);
    end
endmodule

module signextender(outR, inR0,select);
   input wire S1, S0;
   input [31:0] inR0;
   output reg [31:0] outR;
   input [2:0] select;
   wire [31:0] out;
   barrel_shifter bs({24'b000000000000000000000000,inR0[7:0]},out,{1'b0,inR0[11:8]});
   always@(select or inR0)
    begin
   //$display("INSHIFT: %b",inR0);
        case(select)
            3'b000 : outR = inR0;
            3'b001 : begin
            outR= inR0[7:0];
            end
            3'b010 : outR= {5'h00000,inR0[11:0]};
            3'b011 : outR={5'h0000000,inR0[3:0]};
            3'b100 : outR={2'h00,inR0[23:0]};

    endcase
    //$display("OUTSHFT: %b",outR);
     //$display("CONDITIONSELECT WAS: %b",select);
     //$display("CONDITIONMUX OUT: %b",outR);
    end
endmodule

//rotator for 32bitshift001

module barrel_shifter(d,out,m);
  input [31:0]d;
  output [31:0]out,q;
  input[4:0]m;
  wire[4:0] c = m*2;
  mux m1(q[0],d,c);
  mux m2(q[1],{d[0],d[31:1]},c);
  mux m3(q[2],{d[1:0],d[31:2]},c);
  mux m4(q[3],{d[2:0],d[31:3]},c);
  mux m5(q[4],{d[3:0],d[31:4]},c);
  mux m6(q[5],{d[4:0],d[31:5]},c);
  mux m7(q[6],{d[5:0],d[31:6]},c);
  mux m8(q[7],{d[6:0],d[31:7]},c);
  mux m9(q[8],{d[7:0],d[31:8]},c);
  mux m10(q[9],{d[8:0],d[31:9]},c);
  mux m11(q[10],{d[9:0],d[31:10]},c);
  mux m12(q[11],{d[10:0],d[31:11]},c);
  mux m13(q[12],{d[11:0],d[31:12]},c);
  mux m14(q[13],{d[12:0],d[31:13]},c);
  mux m15(q[14],{d[13:0],d[31:14]},c);
  mux m16(q[15],{d[14:0],d[31:15]},c);
  mux m17(q[16],{d[15:0],d[31:16]},c);
  mux m18(q[17],{d[16:0],d[31:17]},c);
  mux m19(q[18],{d[17:0],d[31:18]},c);
  mux m20(q[19],{d[18:0],d[31:19]},c);
  mux m21(q[20],{d[19:0],d[31:20]},c);
  mux m22(q[21],{d[20:0],d[31:21]},c);
  mux m23(q[22],{d[21:0],d[31:22]},c);
  mux m24(q[23],{d[22:0],d[31:23]},c);
  mux m25(q[24],{d[23:0],d[31:24]},c);
  mux m26(q[25],{d[24:0],d[31:25]},c);
  mux m27(q[26],{d[25:0],d[31:26]},c);
  mux m28(q[27],{d[26:0],d[31:27]},c);
  mux m29(q[28],{d[27:0],d[31:28]},c);
  mux m30(q[29],{d[28:0],d[31:29]},c);
  mux m31(q[30],{d[29:0],d[31:30]},c);
  mux m32(q[31],{d[30:0],d[31:31]},c);


  assign out=q;
  always@(out)
  begin
  //$display("BARR: %b",out);
  end
endmodule

module mux(y,d,c);
  input[31:0]d;
  output y;
  reg y;
  input [4:0]c;
  always @ (c)
  begin
    if (c==5'b00000)
      y = d[0];
    else if (c==5'b00001)
      y = d[1];
      else if (c==5'b00010)
      y = d[2];
      else if (c==5'b00011)
      y = d[3];
      else if (c==5'b00100)
      y = d[4];
      else if (c==5'b00101)
      y = d[5];
      else if (c==5'b00110)
      y = d[6];
      else if (c==5'b00111)
      y = d[7];
      else if (c==5'b01000)
      y = d[8];
      else if (c==5'b01001)
      y = d[9];
      else if (c==5'b01010)
      y = d[10];
      else if (c==5'b01011)
      y = d[11];
      else if (c==5'b01100)
      y = d[12];
      else if (c==5'b01101)
      y = d[13];
      else if (c==5'b01110)
      y = d[14];
      else if (c==5'b01111)
      y = d[15];
      else if (c==5'b10000)
      y = d[16];
      else if (c==5'b10001)
      y = d[17];
      else if (c==5'b10010)
      y = d[18];
      else if (c==5'b10011)
      y = d[19];
      else if (c==5'b10100)
      y = d[20];
      else if (c==5'b10101)
      y = d[21];
      else if (c==5'b10110)
      y = d[22];
      else if (c==5'b10111)
      y = d[23];
      else if (c==5'b11000)
      y = d[24];
      else if (c==5'b11001)
      y = d[25];
      else if (c==5'b11010)
      y = d[26];
      else if (c==5'b11011)
      y = d[27];
      else if (c==5'b11100)
      y = d[28];
      else if (c==5'b11101)
      y = d[29];
      else if (c==5'b11110)
      y = d[30];
      else if (c==5'b11111)
      y = d[31];

    end
  endmodule

module instructionRegister(in,out,IREn,clk);
input [31:0] in;
output reg [31:0] out;
input wire IREn,clk;
always@(posedge clk)
begin
if(IREn==1'b1 && in!=32'b00000000000000000000000000001011 && in!=32'b00001011000001010000010000000100)
begin
//$display("INSTRUCTION: %b",iDATAn);
 out = in;
 end
 end
endmodule

module MAR(in,out,enable);
input [31:0] in;
input wire enable;
output reg [7:0] out;
always@(in)
begin
if(enable==1'b1)
begin

//$display("MAR: %d",in[7:0]);
 out = in[7:0];
 end
 end
endmodule

module main;
  wire [7:0] state;
  wire [7:0] stateEncoder;
  wire [31:0] instruction;
  wire [31:0] out;
  wire [7:0] outMux;
  wire MBS,MUXMDR,MDREn,MAREn,IREn,ShiftEn,RFEn,RW,MemEn,MOC, Inv, N2, N1, N0, S1, S0, Sts,iBit, inv, cOutMux,invOut;
  wire [1:0]SignExtSel,MA,MB,MBSMRF;
  wire [2:0] MC;
  wire [1:0] SHF_S;
  wire [5:0] CR;
  wire [4:0] OP;
  wire [7:0] outAdd;
  wire [1:0] M,dataType;
  reg clk, c0, c1;
  //alu+rf
  wire [31:0] portA,portB;
  wire [7:0]currentState;

  //MEMORIA
  wire [31:0]memIn;
  wire [31:0] memOut;
  wire R_W,MOV;
  wire [7:0] address;

  ram_256 ram(memOut,MOC,out,RW,MemEn,address,dataType,stateEncoder);
  MAR mar(out,address,MAREn);
  //Cin
  reg Cin;
  //output
  //Condition codes
  wire zero, n, c, v,R0e,R1e;
  //alu+rfo
  wire [3:0] outMC,outMA;
  wire [31:0] signExtenderOut,R3,R0,R1,R2,R15,outMB,R5;

  instructionRegister ir(memOut,instruction,IREn,clk);
  encoder enc(instruction, stateEncoder);
  conditionMux cMux(cOutMux,1'b0,1'b1,1'b0,1'b0,{S1,S0});
  inverter invert(cOutMux,Inv, invOut);
  nextStAddSel next(M, invOut, N2, N1, N0);
  multiplexer4x1 mux(outMux, stateEncoder, 8'b00000000, CR, outAdd, M);
  multiplexerB b(outMB, portB, signExtenderOut, 32'h00000000, memOut, MB);
  adder add(outMux, 8'b00000001,outAdd);
  ROM rom(R15,R3,zero,dataType,currentState,MA,MB,MC,MBS,MBSMRF,MUXMDR,MDREn,MAREn,IREn,SHF_S,ShiftEn,RFEn,RW,MemEn,MOV, Inv, N2, N1, N0,SignExtSel,CR,OP, outMux,clk,S1,S0,instruction);
  signextender se(signExtenderOut,instruction,SHF_S);
  arithmetic_logic_unit alu(out, zero, n, c, v, portA, outMB, OP, Cin);
  rfMux mc(outMC, instruction[15:12], 4'b1111, instruction[19:16], 4'b1110, MC[1], MC[0]);
  rfMux ma(outMA, instruction[19:16],instruction[15:12], 4'b1111,4'b0000, MA[1], MA[0]);
  registerfile rf(R5,R0,R3,R2,R1,R15,R0e,R1e,out, portA, portB, outMC[3],outMC[2], outMC[1], outMC[0], outMA[3], outMA[2], outMA[1],outMA[0], instruction[3], instruction[2], instruction[1], instruction[0], RFEn, clk);

  initial
  begin
       $display("STATE   |       MAR      |		R15");
       $monitor("%d            %d	%b",currentState,address,R15);
     // $display("R0   |      R1     |    R2      |       R3      |      IR");
     // $monitor("%b            %b        %b      %b          %b",R0,R1,R2,R3,instruction);
     //$display("R2      |       R3       |STATE");
     // $monitor("%b            %b          %d",R2,R3,currentState);
       clk = 0;
        repeat(310)
        begin
            #50 clk = ~clk;
        end
      end
 endmodule
